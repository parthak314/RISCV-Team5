module top (
    input logic clk,
    input logic rst,
    input logic trigger,
    output logic [31:0] a0
);

endmodule