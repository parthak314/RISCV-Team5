module top #(
    parameter DATA_WIDTH = 32
)(
    input logic                     clk,
    input logic                     rst,
    input logic                     trigger,
    output logic [DATA_WIDTH-1:0]   a0
);

endmodule
